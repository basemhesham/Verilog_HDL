`timescale 1ns / 1ps

module seven_segment_decoder(
    input [2:0] inp,
    output reg  seg_a , seg_b , seg_c , seg_d , seg_e , seg_f , seg_g 
);

always @(*) begin
    case (inp)
        3'b000: {seg_a,seg_b,seg_c,seg_d,seg_e,seg_f,seg_g} = 7'b1111110; // 0
        3'b001: {seg_a,seg_b,seg_c,seg_d,seg_e,seg_f,seg_g} = 7'b0110000; // 1
        3'b010: {seg_a,seg_b,seg_c,seg_d,seg_e,seg_f,seg_g} = 7'b1101101; // 2
        3'b011: {seg_a,seg_b,seg_c,seg_d,seg_e,seg_f,seg_g} = 7'b1111001; // 3
        default: 
        {seg_a,seg_b,seg_c,seg_d,seg_e,seg_f,seg_g} = 7'b1001111; // All other values display E
    endcase
end

endmodule

